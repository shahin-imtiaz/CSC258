module try(out);
	output [3:0] out;
	assign out = {2'd10};
endmodule
