module airplane_top (
		CLOCK50,
		VGA_CLK,   						//	VGA Clock
		VGA_HS,							//	VGA H_SYNC
		VGA_VS,							//	VGA V_SYNC
		VGA_BLANK_N,						//	VGA BLANK
		VGA_SYNC_N,						//	VGA SYNC
		VGA_R,   						//	VGA Red[9:0]
		VGA_G,	 						//	VGA Green[9:0]
		VGA_B   						//	VGA Blue[9:0])

		);
		
endmodule





module airplane(clk, reset_n, up, down);
	input CLOCK50;
	input [] KEY;
	
	

endmodule




module datapath(clk, enable, draw, ld_x, ld_y, ld_color, );


endmodule


