module fulladder(a, b, c_in, c_out, s);
	input a;
	input b;
	input c_in;
	output c_out;
	
	assign s = c_in ^ a;
	assign c_out = 
endmodule
