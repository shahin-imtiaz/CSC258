module try(out);
	output [25:0] out;
	assign out = 26'd49999999;
endmodule
