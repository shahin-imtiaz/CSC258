module airplane(clk, reset_n, up, down);
	input CLOCK50;
	input [] KEY;
	
	

endmodule
